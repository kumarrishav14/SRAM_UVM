`include "uvm_macros.svh"
`include "sram_intf.sv"
`include "slave.sv"
`include "sram_trans.sv"
`include "sram_sequence.sv"
`include "sram_driver.sv"
`include "sram_monitor.sv"
`include "sram_agent.sv"
`include "sram_rm.sv"
`include "sram_scb.sv"
`include "sram_fc.sv"
`include "sram_env.sv"
`include "sram_test.sv"